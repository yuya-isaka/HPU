
`default_nettype none


module pop_count
    #(

         // ハイパーベクトルの次元数
         parameter DIM = 1023

     )
     (

         // in
         input wire                     clk,
         input wire                     exec,
         input wire [ DIM:0 ]           data,

         // out
         output wire [ 10:0 ]          result

     );


    reg [ 2:0] stage_1_1;
    reg [ 2:0] stage_1_2;
    reg [ 2:0] stage_1_3;
    reg [ 2:0] stage_1_4;
    reg [ 2:0] stage_1_5;
    reg [ 2:0] stage_1_6;
    reg [ 2:0] stage_1_7;
    reg [ 2:0] stage_1_8;
    reg [ 2:0] stage_1_9;
    reg [ 2:0] stage_1_10;
    reg [ 2:0] stage_1_11;
    reg [ 2:0] stage_1_12;
    reg [ 2:0] stage_1_13;
    reg [ 2:0] stage_1_14;
    reg [ 2:0] stage_1_15;
    reg [ 2:0] stage_1_16;
    reg [ 2:0] stage_1_17;
    reg [ 2:0] stage_1_18;
    reg [ 2:0] stage_1_19;
    reg [ 2:0] stage_1_20;
    reg [ 2:0] stage_1_21;
    reg [ 2:0] stage_1_22;
    reg [ 2:0] stage_1_23;
    reg [ 2:0] stage_1_24;
    reg [ 2:0] stage_1_25;
    reg [ 2:0] stage_1_26;
    reg [ 2:0] stage_1_27;
    reg [ 2:0] stage_1_28;
    reg [ 2:0] stage_1_29;
    reg [ 2:0] stage_1_30;
    reg [ 2:0] stage_1_31;
    reg [ 2:0] stage_1_32;
    reg [ 2:0] stage_1_33;
    reg [ 2:0] stage_1_34;
    reg [ 2:0] stage_1_35;
    reg [ 2:0] stage_1_36;
    reg [ 2:0] stage_1_37;
    reg [ 2:0] stage_1_38;
    reg [ 2:0] stage_1_39;
    reg [ 2:0] stage_1_40;
    reg [ 2:0] stage_1_41;
    reg [ 2:0] stage_1_42;
    reg [ 2:0] stage_1_43;
    reg [ 2:0] stage_1_44;
    reg [ 2:0] stage_1_45;
    reg [ 2:0] stage_1_46;
    reg [ 2:0] stage_1_47;
    reg [ 2:0] stage_1_48;
    reg [ 2:0] stage_1_49;
    reg [ 2:0] stage_1_50;
    reg [ 2:0] stage_1_51;
    reg [ 2:0] stage_1_52;
    reg [ 2:0] stage_1_53;
    reg [ 2:0] stage_1_54;
    reg [ 2:0] stage_1_55;
    reg [ 2:0] stage_1_56;
    reg [ 2:0] stage_1_57;
    reg [ 2:0] stage_1_58;
    reg [ 2:0] stage_1_59;
    reg [ 2:0] stage_1_60;
    reg [ 2:0] stage_1_61;
    reg [ 2:0] stage_1_62;
    reg [ 2:0] stage_1_63;
    reg [ 2:0] stage_1_64;
    reg [ 2:0] stage_1_65;
    reg [ 2:0] stage_1_66;
    reg [ 2:0] stage_1_67;
    reg [ 2:0] stage_1_68;
    reg [ 2:0] stage_1_69;
    reg [ 2:0] stage_1_70;
    reg [ 2:0] stage_1_71;
    reg [ 2:0] stage_1_72;
    reg [ 2:0] stage_1_73;
    reg [ 2:0] stage_1_74;
    reg [ 2:0] stage_1_75;
    reg [ 2:0] stage_1_76;
    reg [ 2:0] stage_1_77;
    reg [ 2:0] stage_1_78;
    reg [ 2:0] stage_1_79;
    reg [ 2:0] stage_1_80;
    reg [ 2:0] stage_1_81;
    reg [ 2:0] stage_1_82;
    reg [ 2:0] stage_1_83;
    reg [ 2:0] stage_1_84;
    reg [ 2:0] stage_1_85;
    reg [ 2:0] stage_1_86;
    reg [ 2:0] stage_1_87;
    reg [ 2:0] stage_1_88;
    reg [ 2:0] stage_1_89;
    reg [ 2:0] stage_1_90;
    reg [ 2:0] stage_1_91;
    reg [ 2:0] stage_1_92;
    reg [ 2:0] stage_1_93;
    reg [ 2:0] stage_1_94;
    reg [ 2:0] stage_1_95;
    reg [ 2:0] stage_1_96;
    reg [ 2:0] stage_1_97;
    reg [ 2:0] stage_1_98;
    reg [ 2:0] stage_1_99;
    reg [ 2:0] stage_1_100;
    reg [ 2:0] stage_1_101;
    reg [ 2:0] stage_1_102;
    reg [ 2:0] stage_1_103;
    reg [ 2:0] stage_1_104;
    reg [ 2:0] stage_1_105;
    reg [ 2:0] stage_1_106;
    reg [ 2:0] stage_1_107;
    reg [ 2:0] stage_1_108;
    reg [ 2:0] stage_1_109;
    reg [ 2:0] stage_1_110;
    reg [ 2:0] stage_1_111;
    reg [ 2:0] stage_1_112;
    reg [ 2:0] stage_1_113;
    reg [ 2:0] stage_1_114;
    reg [ 2:0] stage_1_115;
    reg [ 2:0] stage_1_116;
    reg [ 2:0] stage_1_117;
    reg [ 2:0] stage_1_118;
    reg [ 2:0] stage_1_119;
    reg [ 2:0] stage_1_120;
    reg [ 2:0] stage_1_121;
    reg [ 2:0] stage_1_122;
    reg [ 2:0] stage_1_123;
    reg [ 2:0] stage_1_124;
    reg [ 2:0] stage_1_125;
    reg [ 2:0] stage_1_126;
    reg [ 2:0] stage_1_127;
    reg [ 2:0] stage_1_128;
    reg [ 2:0] stage_1_129;
    reg [ 2:0] stage_1_130;
    reg [ 2:0] stage_1_131;
    reg [ 2:0] stage_1_132;
    reg [ 2:0] stage_1_133;
    reg [ 2:0] stage_1_134;
    reg [ 2:0] stage_1_135;
    reg [ 2:0] stage_1_136;
    reg [ 2:0] stage_1_137;
    reg [ 2:0] stage_1_138;
    reg [ 2:0] stage_1_139;
    reg [ 2:0] stage_1_140;
    reg [ 2:0] stage_1_141;
    reg [ 2:0] stage_1_142;
    reg [ 2:0] stage_1_143;
    reg [ 2:0] stage_1_144;
    reg [ 2:0] stage_1_145;
    reg [ 2:0] stage_1_146;
    reg [ 2:0] stage_1_147;
    reg [ 2:0] stage_1_148;
    reg [ 2:0] stage_1_149;
    reg [ 2:0] stage_1_150;
    reg [ 2:0] stage_1_151;
    reg [ 2:0] stage_1_152;
    reg [ 2:0] stage_1_153;
    reg [ 2:0] stage_1_154;
    reg [ 2:0] stage_1_155;
    reg [ 2:0] stage_1_156;
    reg [ 2:0] stage_1_157;
    reg [ 2:0] stage_1_158;
    reg [ 2:0] stage_1_159;
    reg [ 2:0] stage_1_160;
    reg [ 2:0] stage_1_161;
    reg [ 2:0] stage_1_162;
    reg [ 2:0] stage_1_163;
    reg [ 2:0] stage_1_164;
    reg [ 2:0] stage_1_165;
    reg [ 2:0] stage_1_166;
    reg [ 2:0] stage_1_167;
    reg [ 2:0] stage_1_168;
    reg [ 2:0] stage_1_169;
    reg [ 2:0] stage_1_170;
    reg [ 2:0] stage_1_171;
    reg [ 2:0] stage_1_172;
    reg [ 2:0] stage_1_173;
    reg [ 2:0] stage_1_174;
    reg [ 2:0] stage_1_175;
    reg [ 2:0] stage_1_176;
    reg [ 2:0] stage_1_177;
    reg [ 2:0] stage_1_178;
    reg [ 2:0] stage_1_179;
    reg [ 2:0] stage_1_180;
    reg [ 2:0] stage_1_181;
    reg [ 2:0] stage_1_182;
    reg [ 2:0] stage_1_183;
    reg [ 2:0] stage_1_184;
    reg [ 2:0] stage_1_185;
    reg [ 2:0] stage_1_186;
    reg [ 2:0] stage_1_187;
    reg [ 2:0] stage_1_188;
    reg [ 2:0] stage_1_189;
    reg [ 2:0] stage_1_190;
    reg [ 2:0] stage_1_191;
    reg [ 2:0] stage_1_192;
    reg [ 2:0] stage_1_193;
    reg [ 2:0] stage_1_194;
    reg [ 2:0] stage_1_195;
    reg [ 2:0] stage_1_196;
    reg [ 2:0] stage_1_197;
    reg [ 2:0] stage_1_198;
    reg [ 2:0] stage_1_199;
    reg [ 2:0] stage_1_200;
    reg [ 2:0] stage_1_201;
    reg [ 2:0] stage_1_202;
    reg [ 2:0] stage_1_203;
    reg [ 2:0] stage_1_204;
    reg [ 2:0] stage_1_205;
    reg [ 2:0] stage_1_206;
    reg [ 2:0] stage_1_207;
    reg [ 2:0] stage_1_208;
    reg [ 2:0] stage_1_209;
    reg [ 2:0] stage_1_210;
    reg [ 2:0] stage_1_211;
    reg [ 2:0] stage_1_212;
    reg [ 2:0] stage_1_213;
    reg [ 2:0] stage_1_214;
    reg [ 2:0] stage_1_215;
    reg [ 2:0] stage_1_216;
    reg [ 2:0] stage_1_217;
    reg [ 2:0] stage_1_218;
    reg [ 2:0] stage_1_219;
    reg [ 2:0] stage_1_220;
    reg [ 2:0] stage_1_221;
    reg [ 2:0] stage_1_222;
    reg [ 2:0] stage_1_223;
    reg [ 2:0] stage_1_224;
    reg [ 2:0] stage_1_225;
    reg [ 2:0] stage_1_226;
    reg [ 2:0] stage_1_227;
    reg [ 2:0] stage_1_228;
    reg [ 2:0] stage_1_229;
    reg [ 2:0] stage_1_230;
    reg [ 2:0] stage_1_231;
    reg [ 2:0] stage_1_232;
    reg [ 2:0] stage_1_233;
    reg [ 2:0] stage_1_234;
    reg [ 2:0] stage_1_235;
    reg [ 2:0] stage_1_236;
    reg [ 2:0] stage_1_237;
    reg [ 2:0] stage_1_238;
    reg [ 2:0] stage_1_239;
    reg [ 2:0] stage_1_240;
    reg [ 2:0] stage_1_241;
    reg [ 2:0] stage_1_242;
    reg [ 2:0] stage_1_243;
    reg [ 2:0] stage_1_244;
    reg [ 2:0] stage_1_245;
    reg [ 2:0] stage_1_246;
    reg [ 2:0] stage_1_247;
    reg [ 2:0] stage_1_248;
    reg [ 2:0] stage_1_249;
    reg [ 2:0] stage_1_250;
    reg [ 2:0] stage_1_251;
    reg [ 2:0] stage_1_252;
    reg [ 2:0] stage_1_253;
    reg [ 2:0] stage_1_254;
    reg [ 2:0] stage_1_255;
    reg [ 2:0] stage_1_256;

    always_ff @( posedge clk ) begin

                  if ( exec) begin
                      stage_1_1 <= data[ 0] + data[ 1] + data[ 2] + data[ 3 ];
                      stage_1_2 <= data[ 4] + data[ 5] + data[ 6] + data[ 7 ];
                      stage_1_3 <= data[ 8] + data[ 9] + data[ 10] + data[ 11 ];
                      stage_1_4 <= data[ 12] + data[ 13] + data[ 14] + data[ 15 ];
                      stage_1_5 <= data[ 16] + data[ 17] + data[ 18] + data[ 19 ];
                      stage_1_6 <= data[ 20] + data[ 21] + data[ 22] + data[ 23 ];
                      stage_1_7 <= data[ 24] + data[ 25] + data[ 26] + data[ 27 ];
                      stage_1_8 <= data[ 28] + data[ 29] + data[ 30] + data[ 31 ];
                      stage_1_9 <= data[ 32] + data[ 33] + data[ 34] + data[ 35 ];
                      stage_1_10 <= data[ 36] + data[ 37] + data[ 38] + data[ 39 ];
                      stage_1_11 <= data[ 40] + data[ 41] + data[ 42] + data[ 43 ];
                      stage_1_12 <= data[ 44] + data[ 45] + data[ 46] + data[ 47 ];
                      stage_1_13 <= data[ 48] + data[ 49] + data[ 50] + data[ 51 ];
                      stage_1_14 <= data[ 52] + data[ 53] + data[ 54] + data[ 55 ];
                      stage_1_15 <= data[ 56] + data[ 57] + data[ 58] + data[ 59 ];
                      stage_1_16 <= data[ 60] + data[ 61] + data[ 62] + data[ 63 ];
                      stage_1_17 <= data[ 64] + data[ 65] + data[ 66] + data[ 67 ];
                      stage_1_18 <= data[ 68] + data[ 69] + data[ 70] + data[ 71 ];
                      stage_1_19 <= data[ 72] + data[ 73] + data[ 74] + data[ 75 ];
                      stage_1_20 <= data[ 76] + data[ 77] + data[ 78] + data[ 79 ];
                      stage_1_21 <= data[ 80] + data[ 81] + data[ 82] + data[ 83 ];
                      stage_1_22 <= data[ 84] + data[ 85] + data[ 86] + data[ 87 ];
                      stage_1_23 <= data[ 88] + data[ 89] + data[ 90] + data[ 91 ];
                      stage_1_24 <= data[ 92] + data[ 93] + data[ 94] + data[ 95 ];
                      stage_1_25 <= data[ 96] + data[ 97] + data[ 98] + data[ 99 ];
                      stage_1_26 <= data[ 100] + data[ 101] + data[ 102] + data[ 103 ];
                      stage_1_27 <= data[ 104] + data[ 105] + data[ 106] + data[ 107 ];
                      stage_1_28 <= data[ 108] + data[ 109] + data[ 110] + data[ 111 ];
                      stage_1_29 <= data[ 112] + data[ 113] + data[ 114] + data[ 115 ];
                      stage_1_30 <= data[ 116] + data[ 117] + data[ 118] + data[ 119 ];
                      stage_1_31 <= data[ 120] + data[ 121] + data[ 122] + data[ 123 ];
                      stage_1_32 <= data[ 124] + data[ 125] + data[ 126] + data[ 127 ];
                      stage_1_33 <= data[ 128] + data[ 129] + data[ 130] + data[ 131 ];
                      stage_1_34 <= data[ 132] + data[ 133] + data[ 134] + data[ 135 ];
                      stage_1_35 <= data[ 136] + data[ 137] + data[ 138] + data[ 139 ];
                      stage_1_36 <= data[ 140] + data[ 141] + data[ 142] + data[ 143 ];
                      stage_1_37 <= data[ 144] + data[ 145] + data[ 146] + data[ 147 ];
                      stage_1_38 <= data[ 148] + data[ 149] + data[ 150] + data[ 151 ];
                      stage_1_39 <= data[ 152] + data[ 153] + data[ 154] + data[ 155 ];
                      stage_1_40 <= data[ 156] + data[ 157] + data[ 158] + data[ 159 ];
                      stage_1_41 <= data[ 160] + data[ 161] + data[ 162] + data[ 163 ];
                      stage_1_42 <= data[ 164] + data[ 165] + data[ 166] + data[ 167 ];
                      stage_1_43 <= data[ 168] + data[ 169] + data[ 170] + data[ 171 ];
                      stage_1_44 <= data[ 172] + data[ 173] + data[ 174] + data[ 175 ];
                      stage_1_45 <= data[ 176] + data[ 177] + data[ 178] + data[ 179 ];
                      stage_1_46 <= data[ 180] + data[ 181] + data[ 182] + data[ 183 ];
                      stage_1_47 <= data[ 184] + data[ 185] + data[ 186] + data[ 187 ];
                      stage_1_48 <= data[ 188] + data[ 189] + data[ 190] + data[ 191 ];
                      stage_1_49 <= data[ 192] + data[ 193] + data[ 194] + data[ 195 ];
                      stage_1_50 <= data[ 196] + data[ 197] + data[ 198] + data[ 199 ];
                      stage_1_51 <= data[ 200] + data[ 201] + data[ 202] + data[ 203 ];
                      stage_1_52 <= data[ 204] + data[ 205] + data[ 206] + data[ 207 ];
                      stage_1_53 <= data[ 208] + data[ 209] + data[ 210] + data[ 211 ];
                      stage_1_54 <= data[ 212] + data[ 213] + data[ 214] + data[ 215 ];
                      stage_1_55 <= data[ 216] + data[ 217] + data[ 218] + data[ 219 ];
                      stage_1_56 <= data[ 220] + data[ 221] + data[ 222] + data[ 223 ];
                      stage_1_57 <= data[ 224] + data[ 225] + data[ 226] + data[ 227 ];
                      stage_1_58 <= data[ 228] + data[ 229] + data[ 230] + data[ 231 ];
                      stage_1_59 <= data[ 232] + data[ 233] + data[ 234] + data[ 235 ];
                      stage_1_60 <= data[ 236] + data[ 237] + data[ 238] + data[ 239 ];
                      stage_1_61 <= data[ 240] + data[ 241] + data[ 242] + data[ 243 ];
                      stage_1_62 <= data[ 244] + data[ 245] + data[ 246] + data[ 247 ];
                      stage_1_63 <= data[ 248] + data[ 249] + data[ 250] + data[ 251 ];
                      stage_1_64 <= data[ 252] + data[ 253] + data[ 254] + data[ 255 ];
                      stage_1_65 <= data[ 256] + data[ 257] + data[ 258] + data[ 259 ];
                      stage_1_66 <= data[ 260] + data[ 261] + data[ 262] + data[ 263 ];
                      stage_1_67 <= data[ 264] + data[ 265] + data[ 266] + data[ 267 ];
                      stage_1_68 <= data[ 268] + data[ 269] + data[ 270] + data[ 271 ];
                      stage_1_69 <= data[ 272] + data[ 273] + data[ 274] + data[ 275 ];
                      stage_1_70 <= data[ 276] + data[ 277] + data[ 278] + data[ 279 ];
                      stage_1_71 <= data[ 280] + data[ 281] + data[ 282] + data[ 283 ];
                      stage_1_72 <= data[ 284] + data[ 285] + data[ 286] + data[ 287 ];
                      stage_1_73 <= data[ 288] + data[ 289] + data[ 290] + data[ 291 ];
                      stage_1_74 <= data[ 292] + data[ 293] + data[ 294] + data[ 295 ];
                      stage_1_75 <= data[ 296] + data[ 297] + data[ 298] + data[ 299 ];
                      stage_1_76 <= data[ 300] + data[ 301] + data[ 302] + data[ 303 ];
                      stage_1_77 <= data[ 304] + data[ 305] + data[ 306] + data[ 307 ];
                      stage_1_78 <= data[ 308] + data[ 309] + data[ 310] + data[ 311 ];
                      stage_1_79 <= data[ 312] + data[ 313] + data[ 314] + data[ 315 ];
                      stage_1_80 <= data[ 316] + data[ 317] + data[ 318] + data[ 319 ];
                      stage_1_81 <= data[ 320] + data[ 321] + data[ 322] + data[ 323 ];
                      stage_1_82 <= data[ 324] + data[ 325] + data[ 326] + data[ 327 ];
                      stage_1_83 <= data[ 328] + data[ 329] + data[ 330] + data[ 331 ];
                      stage_1_84 <= data[ 332] + data[ 333] + data[ 334] + data[ 335 ];
                      stage_1_85 <= data[ 336] + data[ 337] + data[ 338] + data[ 339 ];
                      stage_1_86 <= data[ 340] + data[ 341] + data[ 342] + data[ 343 ];
                      stage_1_87 <= data[ 344] + data[ 345] + data[ 346] + data[ 347 ];
                      stage_1_88 <= data[ 348] + data[ 349] + data[ 350] + data[ 351 ];
                      stage_1_89 <= data[ 352] + data[ 353] + data[ 354] + data[ 355 ];
                      stage_1_90 <= data[ 356] + data[ 357] + data[ 358] + data[ 359 ];
                      stage_1_91 <= data[ 360] + data[ 361] + data[ 362] + data[ 363 ];
                      stage_1_92 <= data[ 364] + data[ 365] + data[ 366] + data[ 367 ];
                      stage_1_93 <= data[ 368] + data[ 369] + data[ 370] + data[ 371 ];
                      stage_1_94 <= data[ 372] + data[ 373] + data[ 374] + data[ 375 ];
                      stage_1_95 <= data[ 376] + data[ 377] + data[ 378] + data[ 379 ];
                      stage_1_96 <= data[ 380] + data[ 381] + data[ 382] + data[ 383 ];
                      stage_1_97 <= data[ 384] + data[ 385] + data[ 386] + data[ 387 ];
                      stage_1_98 <= data[ 388] + data[ 389] + data[ 390] + data[ 391 ];
                      stage_1_99 <= data[ 392] + data[ 393] + data[ 394] + data[ 395 ];
                      stage_1_100 <= data[ 396] + data[ 397] + data[ 398] + data[ 399 ];
                      stage_1_101 <= data[ 400] + data[ 401] + data[ 402] + data[ 403 ];
                      stage_1_102 <= data[ 404] + data[ 405] + data[ 406] + data[ 407 ];
                      stage_1_103 <= data[ 408] + data[ 409] + data[ 410] + data[ 411 ];
                      stage_1_104 <= data[ 412] + data[ 413] + data[ 414] + data[ 415 ];
                      stage_1_105 <= data[ 416] + data[ 417] + data[ 418] + data[ 419 ];
                      stage_1_106 <= data[ 420] + data[ 421] + data[ 422] + data[ 423 ];
                      stage_1_107 <= data[ 424] + data[ 425] + data[ 426] + data[ 427 ];
                      stage_1_108 <= data[ 428] + data[ 429] + data[ 430] + data[ 431 ];
                      stage_1_109 <= data[ 432] + data[ 433] + data[ 434] + data[ 435 ];
                      stage_1_110 <= data[ 436] + data[ 437] + data[ 438] + data[ 439 ];
                      stage_1_111 <= data[ 440] + data[ 441] + data[ 442] + data[ 443 ];
                      stage_1_112 <= data[ 444] + data[ 445] + data[ 446] + data[ 447 ];
                      stage_1_113 <= data[ 448] + data[ 449] + data[ 450] + data[ 451 ];
                      stage_1_114 <= data[ 452] + data[ 453] + data[ 454] + data[ 455 ];
                      stage_1_115 <= data[ 456] + data[ 457] + data[ 458] + data[ 459 ];
                      stage_1_116 <= data[ 460] + data[ 461] + data[ 462] + data[ 463 ];
                      stage_1_117 <= data[ 464] + data[ 465] + data[ 466] + data[ 467 ];
                      stage_1_118 <= data[ 468] + data[ 469] + data[ 470] + data[ 471 ];
                      stage_1_119 <= data[ 472] + data[ 473] + data[ 474] + data[ 475 ];
                      stage_1_120 <= data[ 476] + data[ 477] + data[ 478] + data[ 479 ];
                      stage_1_121 <= data[ 480] + data[ 481] + data[ 482] + data[ 483 ];
                      stage_1_122 <= data[ 484] + data[ 485] + data[ 486] + data[ 487 ];
                      stage_1_123 <= data[ 488] + data[ 489] + data[ 490] + data[ 491 ];
                      stage_1_124 <= data[ 492] + data[ 493] + data[ 494] + data[ 495 ];
                      stage_1_125 <= data[ 496] + data[ 497] + data[ 498] + data[ 499 ];
                      stage_1_126 <= data[ 500] + data[ 501] + data[ 502] + data[ 503 ];
                      stage_1_127 <= data[ 504] + data[ 505] + data[ 506] + data[ 507 ];
                      stage_1_128 <= data[ 508] + data[ 509] + data[ 510] + data[ 511 ];
                      stage_1_129 <= data[ 512] + data[ 513] + data[ 514] + data[ 515 ];
                      stage_1_130 <= data[ 516] + data[ 517] + data[ 518] + data[ 519 ];
                      stage_1_131 <= data[ 520] + data[ 521] + data[ 522] + data[ 523 ];
                      stage_1_132 <= data[ 524] + data[ 525] + data[ 526] + data[ 527 ];
                      stage_1_133 <= data[ 528] + data[ 529] + data[ 530] + data[ 531 ];
                      stage_1_134 <= data[ 532] + data[ 533] + data[ 534] + data[ 535 ];
                      stage_1_135 <= data[ 536] + data[ 537] + data[ 538] + data[ 539 ];
                      stage_1_136 <= data[ 540] + data[ 541] + data[ 542] + data[ 543 ];
                      stage_1_137 <= data[ 544] + data[ 545] + data[ 546] + data[ 547 ];
                      stage_1_138 <= data[ 548] + data[ 549] + data[ 550] + data[ 551 ];
                      stage_1_139 <= data[ 552] + data[ 553] + data[ 554] + data[ 555 ];
                      stage_1_140 <= data[ 556] + data[ 557] + data[ 558] + data[ 559 ];
                      stage_1_141 <= data[ 560] + data[ 561] + data[ 562] + data[ 563 ];
                      stage_1_142 <= data[ 564] + data[ 565] + data[ 566] + data[ 567 ];
                      stage_1_143 <= data[ 568] + data[ 569] + data[ 570] + data[ 571 ];
                      stage_1_144 <= data[ 572] + data[ 573] + data[ 574] + data[ 575 ];
                      stage_1_145 <= data[ 576] + data[ 577] + data[ 578] + data[ 579 ];
                      stage_1_146 <= data[ 580] + data[ 581] + data[ 582] + data[ 583 ];
                      stage_1_147 <= data[ 584] + data[ 585] + data[ 586] + data[ 587 ];
                      stage_1_148 <= data[ 588] + data[ 589] + data[ 590] + data[ 591 ];
                      stage_1_149 <= data[ 592] + data[ 593] + data[ 594] + data[ 595 ];
                      stage_1_150 <= data[ 596] + data[ 597] + data[ 598] + data[ 599 ];
                      stage_1_151 <= data[ 600] + data[ 601] + data[ 602] + data[ 603 ];
                      stage_1_152 <= data[ 604] + data[ 605] + data[ 606] + data[ 607 ];
                      stage_1_153 <= data[ 608] + data[ 609] + data[ 610] + data[ 611 ];
                      stage_1_154 <= data[ 612] + data[ 613] + data[ 614] + data[ 615 ];
                      stage_1_155 <= data[ 616] + data[ 617] + data[ 618] + data[ 619 ];
                      stage_1_156 <= data[ 620] + data[ 621] + data[ 622] + data[ 623 ];
                      stage_1_157 <= data[ 624] + data[ 625] + data[ 626] + data[ 627 ];
                      stage_1_158 <= data[ 628] + data[ 629] + data[ 630] + data[ 631 ];
                      stage_1_159 <= data[ 632] + data[ 633] + data[ 634] + data[ 635 ];
                      stage_1_160 <= data[ 636] + data[ 637] + data[ 638] + data[ 639 ];
                      stage_1_161 <= data[ 640] + data[ 641] + data[ 642] + data[ 643 ];
                      stage_1_162 <= data[ 644] + data[ 645] + data[ 646] + data[ 647 ];
                      stage_1_163 <= data[ 648] + data[ 649] + data[ 650] + data[ 651 ];
                      stage_1_164 <= data[ 652] + data[ 653] + data[ 654] + data[ 655 ];
                      stage_1_165 <= data[ 656] + data[ 657] + data[ 658] + data[ 659 ];
                      stage_1_166 <= data[ 660] + data[ 661] + data[ 662] + data[ 663 ];
                      stage_1_167 <= data[ 664] + data[ 665] + data[ 666] + data[ 667 ];
                      stage_1_168 <= data[ 668] + data[ 669] + data[ 670] + data[ 671 ];
                      stage_1_169 <= data[ 672] + data[ 673] + data[ 674] + data[ 675 ];
                      stage_1_170 <= data[ 676] + data[ 677] + data[ 678] + data[ 679 ];
                      stage_1_171 <= data[ 680] + data[ 681] + data[ 682] + data[ 683 ];
                      stage_1_172 <= data[ 684] + data[ 685] + data[ 686] + data[ 687 ];
                      stage_1_173 <= data[ 688] + data[ 689] + data[ 690] + data[ 691 ];
                      stage_1_174 <= data[ 692] + data[ 693] + data[ 694] + data[ 695 ];
                      stage_1_175 <= data[ 696] + data[ 697] + data[ 698] + data[ 699 ];
                      stage_1_176 <= data[ 700] + data[ 701] + data[ 702] + data[ 703 ];
                      stage_1_177 <= data[ 704] + data[ 705] + data[ 706] + data[ 707 ];
                      stage_1_178 <= data[ 708] + data[ 709] + data[ 710] + data[ 711 ];
                      stage_1_179 <= data[ 712] + data[ 713] + data[ 714] + data[ 715 ];
                      stage_1_180 <= data[ 716] + data[ 717] + data[ 718] + data[ 719 ];
                      stage_1_181 <= data[ 720] + data[ 721] + data[ 722] + data[ 723 ];
                      stage_1_182 <= data[ 724] + data[ 725] + data[ 726] + data[ 727 ];
                      stage_1_183 <= data[ 728] + data[ 729] + data[ 730] + data[ 731 ];
                      stage_1_184 <= data[ 732] + data[ 733] + data[ 734] + data[ 735 ];
                      stage_1_185 <= data[ 736] + data[ 737] + data[ 738] + data[ 739 ];
                      stage_1_186 <= data[ 740] + data[ 741] + data[ 742] + data[ 743 ];
                      stage_1_187 <= data[ 744] + data[ 745] + data[ 746] + data[ 747 ];
                      stage_1_188 <= data[ 748] + data[ 749] + data[ 750] + data[ 751 ];
                      stage_1_189 <= data[ 752] + data[ 753] + data[ 754] + data[ 755 ];
                      stage_1_190 <= data[ 756] + data[ 757] + data[ 758] + data[ 759 ];
                      stage_1_191 <= data[ 760] + data[ 761] + data[ 762] + data[ 763 ];
                      stage_1_192 <= data[ 764] + data[ 765] + data[ 766] + data[ 767 ];
                      stage_1_193 <= data[ 768] + data[ 769] + data[ 770] + data[ 771 ];
                      stage_1_194 <= data[ 772] + data[ 773] + data[ 774] + data[ 775 ];
                      stage_1_195 <= data[ 776] + data[ 777] + data[ 778] + data[ 779 ];
                      stage_1_196 <= data[ 780] + data[ 781] + data[ 782] + data[ 783 ];
                      stage_1_197 <= data[ 784] + data[ 785] + data[ 786] + data[ 787 ];
                      stage_1_198 <= data[ 788] + data[ 789] + data[ 790] + data[ 791 ];
                      stage_1_199 <= data[ 792] + data[ 793] + data[ 794] + data[ 795 ];
                      stage_1_200 <= data[ 796] + data[ 797] + data[ 798] + data[ 799 ];
                      stage_1_201 <= data[ 800] + data[ 801] + data[ 802] + data[ 803 ];
                      stage_1_202 <= data[ 804] + data[ 805] + data[ 806] + data[ 807 ];
                      stage_1_203 <= data[ 808] + data[ 809] + data[ 810] + data[ 811 ];
                      stage_1_204 <= data[ 812] + data[ 813] + data[ 814] + data[ 815 ];
                      stage_1_205 <= data[ 816] + data[ 817] + data[ 818] + data[ 819 ];
                      stage_1_206 <= data[ 820] + data[ 821] + data[ 822] + data[ 823 ];
                      stage_1_207 <= data[ 824] + data[ 825] + data[ 826] + data[ 827 ];
                      stage_1_208 <= data[ 828] + data[ 829] + data[ 830] + data[ 831 ];
                      stage_1_209 <= data[ 832] + data[ 833] + data[ 834] + data[ 835 ];
                      stage_1_210 <= data[ 836] + data[ 837] + data[ 838] + data[ 839 ];
                      stage_1_211 <= data[ 840] + data[ 841] + data[ 842] + data[ 843 ];
                      stage_1_212 <= data[ 844] + data[ 845] + data[ 846] + data[ 847 ];
                      stage_1_213 <= data[ 848] + data[ 849] + data[ 850] + data[ 851 ];
                      stage_1_214 <= data[ 852] + data[ 853] + data[ 854] + data[ 855 ];
                      stage_1_215 <= data[ 856] + data[ 857] + data[ 858] + data[ 859 ];
                      stage_1_216 <= data[ 860] + data[ 861] + data[ 862] + data[ 863 ];
                      stage_1_217 <= data[ 864] + data[ 865] + data[ 866] + data[ 867 ];
                      stage_1_218 <= data[ 868] + data[ 869] + data[ 870] + data[ 871 ];
                      stage_1_219 <= data[ 872] + data[ 873] + data[ 874] + data[ 875 ];
                      stage_1_220 <= data[ 876] + data[ 877] + data[ 878] + data[ 879 ];
                      stage_1_221 <= data[ 880] + data[ 881] + data[ 882] + data[ 883 ];
                      stage_1_222 <= data[ 884] + data[ 885] + data[ 886] + data[ 887 ];
                      stage_1_223 <= data[ 888] + data[ 889] + data[ 890] + data[ 891 ];
                      stage_1_224 <= data[ 892] + data[ 893] + data[ 894] + data[ 895 ];
                      stage_1_225 <= data[ 896] + data[ 897] + data[ 898] + data[ 899 ];
                      stage_1_226 <= data[ 900] + data[ 901] + data[ 902] + data[ 903 ];
                      stage_1_227 <= data[ 904] + data[ 905] + data[ 906] + data[ 907 ];
                      stage_1_228 <= data[ 908] + data[ 909] + data[ 910] + data[ 911 ];
                      stage_1_229 <= data[ 912] + data[ 913] + data[ 914] + data[ 915 ];
                      stage_1_230 <= data[ 916] + data[ 917] + data[ 918] + data[ 919 ];
                      stage_1_231 <= data[ 920] + data[ 921] + data[ 922] + data[ 923 ];
                      stage_1_232 <= data[ 924] + data[ 925] + data[ 926] + data[ 927 ];
                      stage_1_233 <= data[ 928] + data[ 929] + data[ 930] + data[ 931 ];
                      stage_1_234 <= data[ 932] + data[ 933] + data[ 934] + data[ 935 ];
                      stage_1_235 <= data[ 936] + data[ 937] + data[ 938] + data[ 939 ];
                      stage_1_236 <= data[ 940] + data[ 941] + data[ 942] + data[ 943 ];
                      stage_1_237 <= data[ 944] + data[ 945] + data[ 946] + data[ 947 ];
                      stage_1_238 <= data[ 948] + data[ 949] + data[ 950] + data[ 951 ];
                      stage_1_239 <= data[ 952] + data[ 953] + data[ 954] + data[ 955 ];
                      stage_1_240 <= data[ 956] + data[ 957] + data[ 958] + data[ 959 ];
                      stage_1_241 <= data[ 960] + data[ 961] + data[ 962] + data[ 963 ];
                      stage_1_242 <= data[ 964] + data[ 965] + data[ 966] + data[ 967 ];
                      stage_1_243 <= data[ 968] + data[ 969] + data[ 970] + data[ 971 ];
                      stage_1_244 <= data[ 972] + data[ 973] + data[ 974] + data[ 975 ];
                      stage_1_245 <= data[ 976] + data[ 977] + data[ 978] + data[ 979 ];
                      stage_1_246 <= data[ 980] + data[ 981] + data[ 982] + data[ 983 ];
                      stage_1_247 <= data[ 984] + data[ 985] + data[ 986] + data[ 987 ];
                      stage_1_248 <= data[ 988] + data[ 989] + data[ 990] + data[ 991 ];
                      stage_1_249 <= data[ 992] + data[ 993] + data[ 994] + data[ 995 ];
                      stage_1_250 <= data[ 996] + data[ 997] + data[ 998] + data[ 999 ];
                      stage_1_251 <= data[ 1000] + data[ 1001] + data[ 1002] + data[ 1003 ];
                      stage_1_252 <= data[ 1004] + data[ 1005] + data[ 1006] + data[ 1007 ];
                      stage_1_253 <= data[ 1008] + data[ 1009] + data[ 1010] + data[ 1011 ];
                      stage_1_254 <= data[ 1012] + data[ 1013] + data[ 1014] + data[ 1015 ];
                      stage_1_255 <= data[ 1016] + data[ 1017] + data[ 1018] + data[ 1019 ];
                      stage_1_256 <= data[ 1020] + data[ 1021] + data[ 1022] + data[ 1023 ];

                  end
              end;

    reg [ 4:0] stage_2_1;
    reg [ 4:0] stage_2_2;
    reg [ 4:0] stage_2_3;
    reg [ 4:0] stage_2_4;
    reg [ 4:0] stage_2_5;
    reg [ 4:0] stage_2_6;
    reg [ 4:0] stage_2_7;
    reg [ 4:0] stage_2_8;
    reg [ 4:0] stage_2_9;
    reg [ 4:0] stage_2_10;
    reg [ 4:0] stage_2_11;
    reg [ 4:0] stage_2_12;
    reg [ 4:0] stage_2_13;
    reg [ 4:0] stage_2_14;
    reg [ 4:0] stage_2_15;
    reg [ 4:0] stage_2_16;
    reg [ 4:0] stage_2_17;
    reg [ 4:0] stage_2_18;
    reg [ 4:0] stage_2_19;
    reg [ 4:0] stage_2_20;
    reg [ 4:0] stage_2_21;
    reg [ 4:0] stage_2_22;
    reg [ 4:0] stage_2_23;
    reg [ 4:0] stage_2_24;
    reg [ 4:0] stage_2_25;
    reg [ 4:0] stage_2_26;
    reg [ 4:0] stage_2_27;
    reg [ 4:0] stage_2_28;
    reg [ 4:0] stage_2_29;
    reg [ 4:0] stage_2_30;
    reg [ 4:0] stage_2_31;
    reg [ 4:0] stage_2_32;
    reg [ 4:0] stage_2_33;
    reg [ 4:0] stage_2_34;
    reg [ 4:0] stage_2_35;
    reg [ 4:0] stage_2_36;
    reg [ 4:0] stage_2_37;
    reg [ 4:0] stage_2_38;
    reg [ 4:0] stage_2_39;
    reg [ 4:0] stage_2_40;
    reg [ 4:0] stage_2_41;
    reg [ 4:0] stage_2_42;
    reg [ 4:0] stage_2_43;
    reg [ 4:0] stage_2_44;
    reg [ 4:0] stage_2_45;
    reg [ 4:0] stage_2_46;
    reg [ 4:0] stage_2_47;
    reg [ 4:0] stage_2_48;
    reg [ 4:0] stage_2_49;
    reg [ 4:0] stage_2_50;
    reg [ 4:0] stage_2_51;
    reg [ 4:0] stage_2_52;
    reg [ 4:0] stage_2_53;
    reg [ 4:0] stage_2_54;
    reg [ 4:0] stage_2_55;
    reg [ 4:0] stage_2_56;
    reg [ 4:0] stage_2_57;
    reg [ 4:0] stage_2_58;
    reg [ 4:0] stage_2_59;
    reg [ 4:0] stage_2_60;
    reg [ 4:0] stage_2_61;
    reg [ 4:0] stage_2_62;
    reg [ 4:0] stage_2_63;
    reg [ 4:0] stage_2_64;

    always_ff @( posedge clk ) begin

                  if ( exec) begin
                      stage_2_1 <= stage_1_1 + stage_1_2 + stage_1_3 + stage_1_4;
                      stage_2_2 <= stage_1_5 + stage_1_6 + stage_1_7 + stage_1_8;
                      stage_2_3 <= stage_1_9 + stage_1_10 + stage_1_11 + stage_1_12;
                      stage_2_4 <= stage_1_13 + stage_1_14 + stage_1_15 + stage_1_16;
                      stage_2_5 <= stage_1_17 + stage_1_18 + stage_1_19 + stage_1_20;
                      stage_2_6 <= stage_1_21 + stage_1_22 + stage_1_23 + stage_1_24;
                      stage_2_7 <= stage_1_25 + stage_1_26 + stage_1_27 + stage_1_28;
                      stage_2_8 <= stage_1_29 + stage_1_30 + stage_1_31 + stage_1_32;
                      stage_2_9 <= stage_1_33 + stage_1_34 + stage_1_35 + stage_1_36;
                      stage_2_10 <= stage_1_37 + stage_1_38 + stage_1_39 + stage_1_40;
                      stage_2_11 <= stage_1_41 + stage_1_42 + stage_1_43 + stage_1_44;
                      stage_2_12 <= stage_1_45 + stage_1_46 + stage_1_47 + stage_1_48;
                      stage_2_13 <= stage_1_49 + stage_1_50 + stage_1_51 + stage_1_52;
                      stage_2_14 <= stage_1_53 + stage_1_54 + stage_1_55 + stage_1_56;
                      stage_2_15 <= stage_1_57 + stage_1_58 + stage_1_59 + stage_1_60;
                      stage_2_16 <= stage_1_61 + stage_1_62 + stage_1_63 + stage_1_64;
                      stage_2_17 <= stage_1_65 + stage_1_66 + stage_1_67 + stage_1_68;
                      stage_2_18 <= stage_1_69 + stage_1_70 + stage_1_71 + stage_1_72;
                      stage_2_19 <= stage_1_73 + stage_1_74 + stage_1_75 + stage_1_76;
                      stage_2_20 <= stage_1_77 + stage_1_78 + stage_1_79 + stage_1_80;
                      stage_2_21 <= stage_1_81 + stage_1_82 + stage_1_83 + stage_1_84;
                      stage_2_22 <= stage_1_85 + stage_1_86 + stage_1_87 + stage_1_88;
                      stage_2_23 <= stage_1_89 + stage_1_90 + stage_1_91 + stage_1_92;
                      stage_2_24 <= stage_1_93 + stage_1_94 + stage_1_95 + stage_1_96;
                      stage_2_25 <= stage_1_97 + stage_1_98 + stage_1_99 + stage_1_100;
                      stage_2_26 <= stage_1_101 + stage_1_102 + stage_1_103 + stage_1_104;
                      stage_2_27 <= stage_1_105 + stage_1_106 + stage_1_107 + stage_1_108;
                      stage_2_28 <= stage_1_109 + stage_1_110 + stage_1_111 + stage_1_112;
                      stage_2_29 <= stage_1_113 + stage_1_114 + stage_1_115 + stage_1_116;
                      stage_2_30 <= stage_1_117 + stage_1_118 + stage_1_119 + stage_1_120;
                      stage_2_31 <= stage_1_121 + stage_1_122 + stage_1_123 + stage_1_124;
                      stage_2_32 <= stage_1_125 + stage_1_126 + stage_1_127 + stage_1_128;
                      stage_2_33 <= stage_1_129 + stage_1_130 + stage_1_131 + stage_1_132;
                      stage_2_34 <= stage_1_133 + stage_1_134 + stage_1_135 + stage_1_136;
                      stage_2_35 <= stage_1_137 + stage_1_138 + stage_1_139 + stage_1_140;
                      stage_2_36 <= stage_1_141 + stage_1_142 + stage_1_143 + stage_1_144;
                      stage_2_37 <= stage_1_145 + stage_1_146 + stage_1_147 + stage_1_148;
                      stage_2_38 <= stage_1_149 + stage_1_150 + stage_1_151 + stage_1_152;
                      stage_2_39 <= stage_1_153 + stage_1_154 + stage_1_155 + stage_1_156;
                      stage_2_40 <= stage_1_157 + stage_1_158 + stage_1_159 + stage_1_160;
                      stage_2_41 <= stage_1_161 + stage_1_162 + stage_1_163 + stage_1_164;
                      stage_2_42 <= stage_1_165 + stage_1_166 + stage_1_167 + stage_1_168;
                      stage_2_43 <= stage_1_169 + stage_1_170 + stage_1_171 + stage_1_172;
                      stage_2_44 <= stage_1_173 + stage_1_174 + stage_1_175 + stage_1_176;
                      stage_2_45 <= stage_1_177 + stage_1_178 + stage_1_179 + stage_1_180;
                      stage_2_46 <= stage_1_181 + stage_1_182 + stage_1_183 + stage_1_184;
                      stage_2_47 <= stage_1_185 + stage_1_186 + stage_1_187 + stage_1_188;
                      stage_2_48 <= stage_1_189 + stage_1_190 + stage_1_191 + stage_1_192;
                      stage_2_49 <= stage_1_193 + stage_1_194 + stage_1_195 + stage_1_196;
                      stage_2_50 <= stage_1_197 + stage_1_198 + stage_1_199 + stage_1_200;
                      stage_2_51 <= stage_1_201 + stage_1_202 + stage_1_203 + stage_1_204;
                      stage_2_52 <= stage_1_205 + stage_1_206 + stage_1_207 + stage_1_208;
                      stage_2_53 <= stage_1_209 + stage_1_210 + stage_1_211 + stage_1_212;
                      stage_2_54 <= stage_1_213 + stage_1_214 + stage_1_215 + stage_1_216;
                      stage_2_55 <= stage_1_217 + stage_1_218 + stage_1_219 + stage_1_220;
                      stage_2_56 <= stage_1_221 + stage_1_222 + stage_1_223 + stage_1_224;
                      stage_2_57 <= stage_1_225 + stage_1_226 + stage_1_227 + stage_1_228;
                      stage_2_58 <= stage_1_229 + stage_1_230 + stage_1_231 + stage_1_232;
                      stage_2_59 <= stage_1_233 + stage_1_234 + stage_1_235 + stage_1_236;
                      stage_2_60 <= stage_1_237 + stage_1_238 + stage_1_239 + stage_1_240;
                      stage_2_61 <= stage_1_241 + stage_1_242 + stage_1_243 + stage_1_244;
                      stage_2_62 <= stage_1_245 + stage_1_246 + stage_1_247 + stage_1_248;
                      stage_2_63 <= stage_1_249 + stage_1_250 + stage_1_251 + stage_1_252;
                      stage_2_64 <= stage_1_253 + stage_1_254 + stage_1_255 + stage_1_256;


                  end
              end;

    reg [ 6:0] stage_3_1;
    reg [ 6:0] stage_3_2;
    reg [ 6:0] stage_3_3;
    reg [ 6:0] stage_3_4;
    reg [ 6:0] stage_3_5;
    reg [ 6:0] stage_3_6;
    reg [ 6:0] stage_3_7;
    reg [ 6:0] stage_3_8;
    reg [ 6:0] stage_3_9;
    reg [ 6:0] stage_3_10;
    reg [ 6:0] stage_3_11;
    reg [ 6:0] stage_3_12;
    reg [ 6:0] stage_3_13;
    reg [ 6:0] stage_3_14;
    reg [ 6:0] stage_3_15;
    reg [ 6:0] stage_3_16;

    always_ff @( posedge clk ) begin

                  if ( exec) begin
                      stage_3_1 <= stage_2_1 + stage_2_2 + stage_2_3 + stage_2_4;
                      stage_3_2 <= stage_2_5 + stage_2_6 + stage_2_7 + stage_2_8;
                      stage_3_3 <= stage_2_9 + stage_2_10 + stage_2_11 + stage_2_12;
                      stage_3_4 <= stage_2_13 + stage_2_14 + stage_2_15 + stage_2_16;
                      stage_3_5 <= stage_2_17 + stage_2_18 + stage_2_19 + stage_2_20;
                      stage_3_6 <= stage_2_21 + stage_2_22 + stage_2_23 + stage_2_24;
                      stage_3_7 <= stage_2_25 + stage_2_26 + stage_2_27 + stage_2_28;
                      stage_3_8 <= stage_2_29 + stage_2_30 + stage_2_31 + stage_2_32;
                      stage_3_9 <= stage_2_33 + stage_2_34 + stage_2_35 + stage_2_36;
                      stage_3_10 <= stage_2_37 + stage_2_38 + stage_2_39 + stage_2_40;
                      stage_3_11 <= stage_2_41 + stage_2_42 + stage_2_43 + stage_2_44;
                      stage_3_12 <= stage_2_45 + stage_2_46 + stage_2_47 + stage_2_48;
                      stage_3_13 <= stage_2_49 + stage_2_50 + stage_2_51 + stage_2_52;
                      stage_3_14 <= stage_2_53 + stage_2_54 + stage_2_55 + stage_2_56;
                      stage_3_15 <= stage_2_57 + stage_2_58 + stage_2_59 + stage_2_60;
                      stage_3_16 <= stage_2_61 + stage_2_62 + stage_2_63 + stage_2_64;
                  end
              end;

    reg [ 8:0] stage_4_1;
    reg [ 8:0] stage_4_2;
    reg [ 8:0] stage_4_3;
    reg [ 8:0] stage_4_4;

    always_ff @( posedge clk ) begin

                  if ( exec) begin
                      stage_4_1 <= stage_3_1 + stage_3_2 + stage_3_3 + stage_3_4;
                      stage_4_2 <= stage_3_5 + stage_3_6 + stage_3_7 + stage_3_8;
                      stage_4_3 <= stage_3_9 + stage_3_10 + stage_3_11 + stage_3_12;
                      stage_4_4 <= stage_3_13 + stage_3_14 + stage_3_15 + stage_3_16;

                  end
              end;

    reg [ 10:0] stage_5_1;

    always_ff @( posedge clk ) begin

                  if ( exec) begin
                      stage_5_1 <= stage_4_1 + stage_4_2 + stage_4_3 + stage_4_4;

                  end
              end;


    assign result = stage_5_1;

endmodule


`default_nettype wire
